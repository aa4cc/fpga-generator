
LIBRARY ieee;
USE ieee.std_logic_1164.all; 
USE ieee.numeric_std.all;

ENTITY Channel IS 
	PORT
	(
		CLK_LOGIC : in std_logic;
		CLK_FREQ  :  in std_logic;
		PHASE_SHIFT_IN : in std_logic_vector(8 downto 0);
		PULSE_WIDTH_IN : in std_logic_vector(8 downto 0);
		RESET : in std_logic;
		OUT_SIGNAL : out std_logic
	);
END Channel;	

architecture arch1 of Channel is

--signal CLK_FREQ : std_logic := '0';


signal phase_shift  : integer range 0 to 360 := 0;
signal duty_width  : integer range 0 to 360 := 180;

signal output : std_logic := '0';

signal newPeriod : std_logic := '0';
signal newPeriodEnable : std_logic := '1';

signal duty_begin : std_logic := '0';
signal duty_on : std_logic := '0';
signal duty_enable : std_logic := '1';


begin


phase_shift <= to_integer(unsigned(PHASE_SHIFT_IN));
duty_width <= to_integer(unsigned(PULSE_WIDTH_IN)) when phase_shift < 361 	else 0;




--OUT_SIGNAL <= output;
OUT_SIGNAL <= duty_on; --and duty_enable;


 shiftPhase : process(CLK_LOGIC, RESET) is
  variable counter : integer range 0 to 400 := 0;
  variable counting : std_logic := '0';
  variable lastFreq : std_logic := '0';
  variable countingLag : std_logic := '0';
  
 
  begin
  
  if reset = '1' then
				--reset
				counter := 0;
				counting := '0';
				lastFreq := '0';
				countingLag := '0';
				duty_begin <= '0';
				duty_enable <= '1';
  else
	  
	  if rising_edge(CLK_LOGIC) then
			if counting = '0' then
				if CLK_FREQ = '1' and lastFreq = '0' then
					if phase_shift = 0 then
						duty_begin <= '1';
					else
						counting := '1';
						counter := phase_shift;
						duty_begin <= '0';
					end if;
					
				else
					counting := '0';
					duty_begin <= '0';
				end if;
			elsif counting = '1' then
				if counter = 1 then
					duty_begin <= '1';
					counting := '0';
				else
					counter := counter - 1;
					duty_begin <= '0';
				end if;
			end if;
	  
	  lastFreq := CLK_FREQ;
	  duty_enable <= not(countingLag);
	  countingLag := counting;
	  --duty_begin <= counting;
			
	  end if;
  end if;
 
  end process shiftPhase;
  
  
  
  
  dutyCycle : process(CLK_LOGIC) is
  variable counter : integer range 0 to 400 := 0;
  variable counting : std_logic := '0';
  variable lastBegin : std_logic := '0';
  variable duty_out : std_logic := '0';
 
  begin
  
  if reset = '1' then
				--reset
				counter := 0;
				counting := '0';
				lastBegin := '0';
				duty_out := '0';
				output <= '0';
				newPeriod <= '0';
				newPeriodEnable <= '1';
				duty_on <= '0';
				duty_enable <= '1';
  else
	  
	  if rising_edge(CLK_LOGIC) then
			if counting = '0' then
				if duty_begin = '1' and lastBegin = '0' then
					if duty_width = 0 then
						--do nothing
					else
						counting := '1';
						counter := duty_width;
						duty_on <= '1';
					end if;
					
				else
					counting := '0';
					duty_on <= '0';
				end if;
			elsif counting = '1' then
				if counter = 1 then
					duty_on <= '0';
					counting := '0';
				else
					counter := counter - 1;
					duty_on <= '1';
				end if;
			end if;
	  
	  lastBegin := duty_begin;
			
	  end if;
  end if;
  end process dutyCycle;
  
  
end arch1;

